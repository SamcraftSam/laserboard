*Photodiode NOISE Analysis Spice Netlist - 2 stages using AD8656

* input signal - photodiode current, and noise source for noise analysis 
IS IN 0 AC 1 PULSE(0 4u 1n 1n 1n 1 2)
VNOISE INP 0 AC 0

VP VCCG 0 2.75
VM VEEG 0 -2.75

* Photodiode model and TIA amplifier circuit 
*Stage 1 
X1 INP IN VCCG VEEG OUT1 AD8656
RSH IN 0 5G
CD IN 0 25p
RF IN OUT1 82.5k
CF IN OUT1 2.7p

*Stage 2 
X2 INP2 INN2 VCCG VEEG OUT AD8656
Rfilt OUT1 INP2 487
Cfilt INP2 0 330p
RF2 OUT INN2 825
RG2 INN2 0 162

* simulation directives 
.NOISE V(OUT) VNOISE DEC 100 10k 105Meg

* AD8656 SPICE Macro-model
* Description: Amplifier
* Generic Desc: 2.7/5V, CMOS, OP, Low Noise, RRIO, 2X
* Developed by: ADSJ HH
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (06/2005)
* Copyright 2010, 2012 by Analog Devices
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement.  Use of this model
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*    
* Parameters modeled include:
*
* END Notes
*
* Node Assignments
*                       noninverting input
*                       |   inverting input
*                       |   |    positive supply
*                       |   |    |   negative supply
*                       |   |    |   |   output
*                       |   |    |   |   |
*                       |   |    |   |   |
.SUBCKT AD8656      	1   2   99  50  45
*
* INPUT STAGE
*
M1  14  7  8  8 PIX L=1E-6 W=1.45E-02
M2  16  2  8  8 PIX L=1E-6 W=1.45E-02
M3  17  7 10 10 NIX L=1E-6 W=1.45E-02
M4  18  2 10 10 NIX L=1E-6 W=1.45E-02
RD1 14 50 8.00E+02
RD2 16 50 8.00E+02
RD3 99 17 8.00E+02
RD4 99 18 8.00E+02
C1  14 16 1.22E-12
C2  17 18 1.22E-12
I1  99  8 5.00E-04
I2  10 50 5.00E-04
V1  99  9 1.141E+00
V2  13 50 1.141E+00
D1   8  9 DX
D2  13 10 DX
EOS  7  1 POLY(4) (22,98) (73,98) (81,98) (70,98) 5.00E-05 1 1 1 1
IOS  1  2 5.00E-13
*
*CMRR=110dB, POLE AT 400 Hz
*
E1  21 98 POLY(2) (1,98) (2,98) 0 3.95E-02 3.95E-02
R10 21 22 3.98E+02
R20 22 98 1.59E-02
C10 21 22 1.00E-06
*
* PSRR=93dB, POLE AT 1500 Hz
*
EPSY 72 98 POLY(1) (99,50) -7.462403795 1.492480759
CPS3 72 73 1.00E-06
RPS3 72 73 1.06E+02
RPS4 73 98 1.59E-03
*
* VOLTAGE NOISE REFERENCE OF 2.7nV/rt(Hz)
*
VN1 80 98 0
RN1 80 98 16.45E-3
HN  81 98 VN1 2.39E+00
RN2 81 98 1
*
* FLICKER NOISE CORNER = 1200 Hz
*
D5  69 98 DNOISE
VSN 69 98 DC 0.6551
H1  70 98 POLY(1) VSN 1.00E-03 1.00E+00
RN  70 98 1
*
* INTERNAL VOLTAGE REFERENCE
*
EREF 98  0 POLY(2) (99,0) (50,0) 0 0.5 0.5
GSY  99 50 POLY(1) (99,50) 1.68E-03 1.10E-06
EVP  97 98 POLY(1) (99,50) 0 0.5
EVN  51 98 POLY(1) (50,99) 0 0.5
*
* GAIN STAGE
*
G1 98 30 POLY(2) (14,16) (17,18) 0 1.68E-04 1.68E-04
R1 30 98 1.00E+06
RZ 30 31 4.58E+01
CF 45 31 1.22E-11
V3 32 30 -4.95E-01
V4 30 33 -1.79E+00
D3 32 97 DX
D4 51 33 DX
*
* OUTPUT STAGE
*
M5  45 46 99 99 POX L=1E-6 W=2.37E-03
M6  45 47 50 50 NOX L=1E-6 W=2.81E-03
EG1 99 46 POLY(1) (98,30) 6.169E-01 1
EG2 47 50 POLY(1) (30,98) 5.934E-01 1
*
* MODELS
*
.MODEL POX PMOS (LEVEL=2,KP=1.00E-05,VTO=-0.328,LAMBDA=0.01,RD=0)
.MODEL NOX NMOS (LEVEL=2,KP=1.00E-05,VTO=+0.328,LAMBDA=0.01,RD=0)
.MODEL PIX PMOS (LEVEL=2,KP=1.00E-05,VTO=-0.5,LAMBDA=0.01)
.MODEL NIX NMOS (LEVEL=2,KP=1.00E-05,VTO=0.5,LAMBDA=0.01)
.MODEL DX D(IS=1E-14,RS=5)
.MODEL DNOISE D(IS=1E-14,RS=0,KF=8.75E-12)
*
*
.ENDS AD8656
*
*




